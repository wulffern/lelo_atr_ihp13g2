magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 3696 2560
use LELOATR_NCH_8CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 1848 480
use LELOATR_NCH_8C1F2 xa2 
transform 1 0 0 0 1 480
box 0 480 1848 1280
use LELOATR_NCH_8C5F0 xa3 
transform 1 0 0 0 1 1280
box 0 1280 1848 2080
use LELOATR_NCH_8CTAPTOP xa4 
transform 1 0 0 0 1 2080
box 0 2080 1848 2560
use LELOATR_NCH_8CTAPBOT xb1 
transform 1 0 1848 0 1 0
box 1848 0 3696 480
use LELOATR_NCH_8C1F2 xb2 
transform 1 0 1848 0 1 480
box 1848 480 3696 1280
use LELOATR_NCH_8C5F0 xb3 
transform 1 0 1848 0 1 1280
box 1848 1280 3696 2080
use LELOATR_NCH_8CTAPTOP xb4 
transform 1 0 1848 0 1 2080
box 1848 2080 3696 2560
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 3696 2560
<< end >>
