magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 3024 2560
use LELOATR_PCH_4CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 1512 480
use LELOATR_PCH_4C1F2 xa2 
transform 1 0 0 0 1 480
box 0 480 1512 1280
use LELOATR_PCH_4C5F0 xa3 
transform 1 0 0 0 1 1280
box 0 1280 1512 2080
use LELOATR_PCH_4CTAPTOP xa4 
transform 1 0 0 0 1 2080
box 0 2080 1512 2560
use LELOATR_PCH_4CTAPBOT xb1 
transform 1 0 1512 0 1 0
box 1512 0 3024 480
use LELOATR_PCH_4C1F2 xb2 
transform 1 0 1512 0 1 480
box 1512 480 3024 1280
use LELOATR_PCH_4C5F0 xb3 
transform 1 0 1512 0 1 1280
box 1512 1280 3024 2080
use LELOATR_PCH_4CTAPTOP xb4 
transform 1 0 1512 0 1 2080
box 1512 2080 3024 2560
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 3024 2560
<< end >>
