magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 1512 800
<< pdiff >>
rect 546 40 966 120
rect 546 120 966 200
rect 546 200 966 280
rect 546 280 966 360
rect 546 360 966 440
rect 546 440 966 520
rect 546 520 966 600
rect 546 600 966 680
rect 546 680 966 760
<< ptap >>
rect -126 -40 126 40
rect 1386 -40 1638 40
rect -126 40 126 120
rect 1386 40 1638 120
rect -126 120 126 200
rect 1386 120 1638 200
rect -126 200 126 280
rect 1386 200 1638 280
rect -126 280 126 360
rect 1386 280 1638 360
rect -126 360 126 440
rect 1386 360 1638 440
rect -126 440 126 520
rect 1386 440 1638 520
rect -126 520 126 600
rect 1386 520 1638 600
rect -126 600 126 680
rect 1386 600 1638 680
rect -126 680 126 760
rect 1386 680 1638 760
rect -126 760 126 840
rect 1386 760 1638 840
<< poly >>
rect 210 140 1302 340
rect 210 460 1302 660
rect 210 -14 1302 14
rect 210 200 294 280
rect 1218 200 1302 280
rect 210 280 294 360
rect 1218 280 1302 360
rect 210 360 294 440
rect 1218 360 1302 440
rect 210 440 294 520
rect 1218 440 1302 520
rect 210 520 294 600
rect 1218 520 1302 600
rect 210 786 1302 814
<< metal2 >>
rect 210 360 294 440
rect 378 600 630 680
rect 882 40 1134 120
rect 210 40 294 120
rect 378 40 630 120
rect 882 40 1134 120
rect 210 120 294 200
rect 378 120 630 200
rect 882 120 1134 200
rect 210 200 294 280
rect 378 200 630 280
rect 882 200 1134 280
rect 210 280 294 360
rect 378 280 630 360
rect 882 280 1134 360
rect 210 360 294 440
rect 378 360 630 440
rect 882 360 1134 440
rect 210 440 294 520
rect 378 440 630 520
rect 882 440 1134 520
rect 210 520 294 600
rect 378 520 630 600
rect 882 520 1134 600
rect 210 600 294 680
rect 378 600 630 680
rect 882 600 1134 680
rect 210 680 294 760
rect 378 680 630 760
rect 882 680 1134 760
<< pc >>
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 1232 300 1288 320
rect 1232 320 1288 340
rect 1232 340 1288 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1232 360 1288 380
rect 1232 380 1288 400
rect 1232 400 1288 420
rect 1232 420 1288 440
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 1232 440 1288 460
rect 1232 460 1288 480
rect 1232 480 1288 500
<< metal1 >>
rect -126 -40 126 40
rect 1386 -40 1638 40
rect -126 40 126 120
rect 378 40 966 120
rect 1386 40 1638 120
rect -126 120 126 200
rect 1386 120 1638 200
rect -126 200 126 280
rect 1386 200 1638 280
rect -126 280 126 360
rect 210 280 294 360
rect 1218 280 1302 360
rect 1386 280 1638 360
rect -126 360 126 440
rect -126 360 126 440
rect 210 360 294 440
rect 546 360 1134 440
rect 1218 360 1302 440
rect 1386 360 1638 440
rect -126 440 126 520
rect 210 440 294 520
rect 1218 440 1302 520
rect 1386 440 1638 520
rect -126 520 126 600
rect 1386 520 1638 600
rect -126 600 126 680
rect 1386 600 1638 680
rect -126 680 126 760
rect 378 680 966 760
rect 1386 680 1638 760
rect -126 760 126 840
rect 1386 760 1638 840
<< ptapc >>
rect -42 200 42 280
rect 1470 200 1554 280
rect -42 280 42 360
rect 1470 280 1554 360
rect -42 360 42 440
rect 1470 360 1554 440
rect -42 440 42 520
rect 1470 440 1554 520
rect -42 520 42 600
rect 1470 520 1554 600
<< ndcontact >>
rect 588 60 630 80
rect 588 80 630 100
rect 630 60 714 80
rect 630 80 714 100
rect 714 60 798 80
rect 714 80 798 100
rect 798 60 882 80
rect 798 80 882 100
rect 882 60 924 80
rect 882 80 924 100
rect 588 380 630 400
rect 588 400 630 420
rect 630 380 714 400
rect 630 400 714 420
rect 714 380 798 400
rect 714 400 798 420
rect 798 380 882 400
rect 798 400 882 420
rect 882 380 924 400
rect 882 400 924 420
rect 588 700 630 720
rect 588 720 630 740
rect 630 700 714 720
rect 630 720 714 740
rect 714 700 798 720
rect 714 720 798 740
rect 798 700 882 720
rect 798 720 882 740
rect 882 700 924 720
rect 882 720 924 740
<< via1 >>
rect 420 48 462 56
rect 420 56 462 64
rect 420 64 462 72
rect 420 72 462 80
rect 420 80 462 88
rect 420 88 462 96
rect 420 96 462 104
rect 420 104 462 112
rect 462 48 546 56
rect 462 56 546 64
rect 462 64 546 72
rect 462 72 546 80
rect 462 80 546 88
rect 462 88 546 96
rect 462 96 546 104
rect 462 104 546 112
rect 546 48 588 56
rect 546 56 588 64
rect 546 64 588 72
rect 546 72 588 80
rect 546 80 588 88
rect 546 88 588 96
rect 546 96 588 104
rect 546 104 588 112
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 924 368 966 376
rect 924 376 966 384
rect 924 384 966 392
rect 924 392 966 400
rect 924 400 966 408
rect 924 408 966 416
rect 924 416 966 424
rect 924 424 966 432
rect 966 368 1050 376
rect 966 376 1050 384
rect 966 384 1050 392
rect 966 392 1050 400
rect 966 400 1050 408
rect 966 408 1050 416
rect 966 416 1050 424
rect 966 424 1050 432
rect 1050 368 1092 376
rect 1050 376 1092 384
rect 1050 384 1092 392
rect 1050 392 1092 400
rect 1050 400 1092 408
rect 1050 408 1092 416
rect 1050 416 1092 424
rect 1050 424 1092 432
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 420 688 462 696
rect 420 696 462 704
rect 420 704 462 712
rect 420 712 462 720
rect 420 720 462 728
rect 420 728 462 736
rect 420 736 462 744
rect 420 744 462 752
rect 462 688 546 696
rect 462 696 546 704
rect 462 704 546 712
rect 462 712 546 720
rect 462 720 546 728
rect 462 728 546 736
rect 462 736 546 744
rect 462 744 546 752
rect 546 688 588 696
rect 546 696 588 704
rect 546 704 588 712
rect 546 712 588 720
rect 546 720 588 728
rect 546 728 588 736
rect 546 736 588 744
rect 546 744 588 752
<< pwell >>
rect -126 -40 1638 840
<< labels >>
flabel metal2 s 210 360 294 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel metal2 s 378 600 630 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel metal1 s -126 360 126 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel metal2 s 882 40 1134 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1512 800
<< end >>
