magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 1848 800
<< pdiff >>
rect 546 200 1302 280
rect 546 280 1302 360
rect 546 360 1302 440
rect 546 440 1302 520
rect 546 520 1302 600
<< ntap >>
rect -126 -40 126 40
rect 1722 -40 1974 40
rect -126 40 126 120
rect 1722 40 1974 120
rect -126 120 126 200
rect 1722 120 1974 200
rect -126 200 126 280
rect 1722 200 1974 280
rect -126 280 126 360
rect 1722 280 1974 360
rect -126 360 126 440
rect 1722 360 1974 440
rect -126 440 126 520
rect 1722 440 1974 520
rect -126 520 126 600
rect 1722 520 1974 600
rect -126 600 126 680
rect 1722 600 1974 680
rect -126 680 126 760
rect 1722 680 1974 760
rect -126 760 126 840
rect 1722 760 1974 840
<< poly >>
rect 210 -14 1638 14
rect 210 146 1638 174
rect 210 306 1638 334
rect 210 466 1638 494
rect 210 626 1638 654
rect 210 786 1638 814
rect 210 280 294 360
rect 1554 280 1638 360
rect 210 360 294 440
rect 1554 360 1638 440
rect 210 440 294 520
rect 1554 440 1638 520
<< metal2 >>
rect 210 360 294 440
rect 378 600 630 680
rect 1218 40 1470 120
rect 210 40 294 120
rect 378 40 630 120
rect 1218 40 1470 120
rect 210 120 294 200
rect 378 120 630 200
rect 1218 120 1470 200
rect 210 200 294 280
rect 378 200 630 280
rect 1218 200 1470 280
rect 210 280 294 360
rect 378 280 630 360
rect 1218 280 1470 360
rect 210 360 294 440
rect 378 360 630 440
rect 1218 360 1470 440
rect 210 440 294 520
rect 378 440 630 520
rect 1218 440 1470 520
rect 210 520 294 600
rect 378 520 630 600
rect 1218 520 1470 600
rect 210 600 294 680
rect 378 600 630 680
rect 1218 600 1470 680
rect 210 680 294 760
rect 378 680 630 760
rect 1218 680 1470 760
<< pc >>
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 1568 300 1624 320
rect 1568 320 1624 340
rect 1568 340 1624 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1568 360 1624 380
rect 1568 380 1624 400
rect 1568 400 1624 420
rect 1568 420 1624 440
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 1568 440 1624 460
rect 1568 460 1624 480
rect 1568 480 1624 500
<< metal1 >>
rect -126 -40 126 40
rect 1722 -40 1974 40
rect -126 40 126 120
rect 1722 40 1974 120
rect -126 120 126 200
rect 1722 120 1974 200
rect -126 200 126 280
rect 378 200 1302 280
rect 1722 200 1974 280
rect -126 280 126 360
rect 210 280 294 360
rect 1554 280 1638 360
rect 1722 280 1974 360
rect -126 360 126 440
rect -126 360 126 440
rect 210 360 294 440
rect 546 360 1470 440
rect 1554 360 1638 440
rect 1722 360 1974 440
rect -126 440 126 520
rect 210 440 294 520
rect 1554 440 1638 520
rect 1722 440 1974 520
rect -126 520 126 600
rect 378 520 1302 600
rect 1722 520 1974 600
rect -126 600 126 680
rect 1722 600 1974 680
rect -126 680 126 760
rect 1722 680 1974 760
rect -126 760 126 840
rect 1722 760 1974 840
<< ntapc >>
rect -42 200 42 280
rect 1806 200 1890 280
rect -42 280 42 360
rect 1806 280 1890 360
rect -42 360 42 440
rect 1806 360 1890 440
rect -42 440 42 520
rect 1806 440 1890 520
rect -42 520 42 600
rect 1806 520 1890 600
<< pdcontact >>
rect 588 220 630 240
rect 588 240 630 260
rect 630 220 714 240
rect 630 240 714 260
rect 714 220 798 240
rect 714 240 798 260
rect 798 220 882 240
rect 798 240 882 260
rect 882 220 966 240
rect 882 240 966 260
rect 966 220 1050 240
rect 966 240 1050 260
rect 1050 220 1134 240
rect 1050 240 1134 260
rect 1134 220 1218 240
rect 1134 240 1218 260
rect 1218 220 1260 240
rect 1218 240 1260 260
rect 588 380 630 400
rect 588 400 630 420
rect 630 380 714 400
rect 630 400 714 420
rect 714 380 798 400
rect 714 400 798 420
rect 798 380 882 400
rect 798 400 882 420
rect 882 380 966 400
rect 882 400 966 420
rect 966 380 1050 400
rect 966 400 1050 420
rect 1050 380 1134 400
rect 1050 400 1134 420
rect 1134 380 1218 400
rect 1134 400 1218 420
rect 1218 380 1260 400
rect 1218 400 1260 420
rect 588 540 630 560
rect 588 560 630 580
rect 630 540 714 560
rect 630 560 714 580
rect 714 540 798 560
rect 714 560 798 580
rect 798 540 882 560
rect 798 560 882 580
rect 882 540 966 560
rect 882 560 966 580
rect 966 540 1050 560
rect 966 560 1050 580
rect 1050 540 1134 560
rect 1050 560 1134 580
rect 1134 540 1218 560
rect 1134 560 1218 580
rect 1218 540 1260 560
rect 1218 560 1260 580
<< via1 >>
rect 420 208 462 216
rect 420 216 462 224
rect 420 224 462 232
rect 420 232 462 240
rect 420 240 462 248
rect 420 248 462 256
rect 420 256 462 264
rect 420 264 462 272
rect 462 208 546 216
rect 462 216 546 224
rect 462 224 546 232
rect 462 232 546 240
rect 462 240 546 248
rect 462 248 546 256
rect 462 256 546 264
rect 462 264 546 272
rect 546 208 588 216
rect 546 216 588 224
rect 546 224 588 232
rect 546 232 588 240
rect 546 240 588 248
rect 546 248 588 256
rect 546 256 588 264
rect 546 264 588 272
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1260 368 1302 376
rect 1260 376 1302 384
rect 1260 384 1302 392
rect 1260 392 1302 400
rect 1260 400 1302 408
rect 1260 408 1302 416
rect 1260 416 1302 424
rect 1260 424 1302 432
rect 1302 368 1386 376
rect 1302 376 1386 384
rect 1302 384 1386 392
rect 1302 392 1386 400
rect 1302 400 1386 408
rect 1302 408 1386 416
rect 1302 416 1386 424
rect 1302 424 1386 432
rect 1386 368 1428 376
rect 1386 376 1428 384
rect 1386 384 1428 392
rect 1386 392 1428 400
rect 1386 400 1428 408
rect 1386 408 1428 416
rect 1386 416 1428 424
rect 1386 424 1428 432
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 420 528 462 536
rect 420 536 462 544
rect 420 544 462 552
rect 420 552 462 560
rect 420 560 462 568
rect 420 568 462 576
rect 420 576 462 584
rect 420 584 462 592
rect 462 528 546 536
rect 462 536 546 544
rect 462 544 546 552
rect 462 552 546 560
rect 462 560 546 568
rect 462 568 546 576
rect 462 576 546 584
rect 462 584 546 592
rect 546 528 588 536
rect 546 536 588 544
rect 546 544 588 552
rect 546 552 588 560
rect 546 560 588 568
rect 546 568 588 576
rect 546 576 588 584
rect 546 584 588 592
<< nwell >>
rect -210 -124 2058 924
<< labels >>
flabel metal2 s 210 360 294 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel metal2 s 378 600 630 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel metal1 s -126 360 126 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel metal2 s 1218 40 1470 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1848 800
<< end >>
