magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 2184 800
<< pdiff >>
rect 546 40 1638 120
rect 546 120 1638 200
rect 546 200 1638 280
rect 546 280 1638 360
rect 546 360 1638 440
rect 546 440 1638 520
rect 546 520 1638 600
rect 546 600 1638 680
rect 546 680 1638 760
<< ptap >>
rect -126 -40 126 40
rect 2058 -40 2310 40
rect -126 40 126 120
rect 2058 40 2310 120
rect -126 120 126 200
rect 2058 120 2310 200
rect -126 200 126 280
rect 2058 200 2310 280
rect -126 280 126 360
rect 2058 280 2310 360
rect -126 360 126 440
rect 2058 360 2310 440
rect -126 440 126 520
rect 2058 440 2310 520
rect -126 520 126 600
rect 2058 520 2310 600
rect -126 600 126 680
rect 2058 600 2310 680
rect -126 680 126 760
rect 2058 680 2310 760
rect -126 760 126 840
rect 2058 760 2310 840
<< poly >>
rect 210 140 1974 340
rect 210 460 1974 660
rect 210 -14 1974 14
rect 210 200 294 280
rect 1890 200 1974 280
rect 210 280 294 360
rect 1890 280 1974 360
rect 210 360 294 440
rect 1890 360 1974 440
rect 210 440 294 520
rect 1890 440 1974 520
rect 210 520 294 600
rect 1890 520 1974 600
rect 210 786 1974 814
<< metal2 >>
rect 210 360 294 440
rect 378 600 630 680
rect 1554 40 1806 120
rect 210 40 294 120
rect 378 40 630 120
rect 1554 40 1806 120
rect 210 120 294 200
rect 378 120 630 200
rect 1554 120 1806 200
rect 210 200 294 280
rect 378 200 630 280
rect 1554 200 1806 280
rect 210 280 294 360
rect 378 280 630 360
rect 1554 280 1806 360
rect 210 360 294 440
rect 378 360 630 440
rect 1554 360 1806 440
rect 210 440 294 520
rect 378 440 630 520
rect 1554 440 1806 520
rect 210 520 294 600
rect 378 520 630 600
rect 1554 520 1806 600
rect 210 600 294 680
rect 378 600 630 680
rect 1554 600 1806 680
rect 210 680 294 760
rect 378 680 630 760
rect 1554 680 1806 760
<< pc >>
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 1904 300 1960 320
rect 1904 320 1960 340
rect 1904 340 1960 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1904 360 1960 380
rect 1904 380 1960 400
rect 1904 400 1960 420
rect 1904 420 1960 440
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 1904 440 1960 460
rect 1904 460 1960 480
rect 1904 480 1960 500
<< metal1 >>
rect -126 -40 126 40
rect 2058 -40 2310 40
rect -126 40 126 120
rect 378 40 1638 120
rect 2058 40 2310 120
rect -126 120 126 200
rect 2058 120 2310 200
rect -126 200 126 280
rect 2058 200 2310 280
rect -126 280 126 360
rect 210 280 294 360
rect 1890 280 1974 360
rect 2058 280 2310 360
rect -126 360 126 440
rect -126 360 126 440
rect 210 360 294 440
rect 546 360 1806 440
rect 1890 360 1974 440
rect 2058 360 2310 440
rect -126 440 126 520
rect 210 440 294 520
rect 1890 440 1974 520
rect 2058 440 2310 520
rect -126 520 126 600
rect 2058 520 2310 600
rect -126 600 126 680
rect 2058 600 2310 680
rect -126 680 126 760
rect 378 680 1638 760
rect 2058 680 2310 760
rect -126 760 126 840
rect 2058 760 2310 840
<< ptapc >>
rect -42 200 42 280
rect 2142 200 2226 280
rect -42 280 42 360
rect 2142 280 2226 360
rect -42 360 42 440
rect 2142 360 2226 440
rect -42 440 42 520
rect 2142 440 2226 520
rect -42 520 42 600
rect 2142 520 2226 600
<< ndcontact >>
rect 588 60 630 80
rect 588 80 630 100
rect 630 60 714 80
rect 630 80 714 100
rect 714 60 798 80
rect 714 80 798 100
rect 798 60 882 80
rect 798 80 882 100
rect 882 60 966 80
rect 882 80 966 100
rect 966 60 1050 80
rect 966 80 1050 100
rect 1050 60 1134 80
rect 1050 80 1134 100
rect 1134 60 1218 80
rect 1134 80 1218 100
rect 1218 60 1302 80
rect 1218 80 1302 100
rect 1302 60 1386 80
rect 1302 80 1386 100
rect 1386 60 1470 80
rect 1386 80 1470 100
rect 1470 60 1554 80
rect 1470 80 1554 100
rect 1554 60 1596 80
rect 1554 80 1596 100
rect 588 380 630 400
rect 588 400 630 420
rect 630 380 714 400
rect 630 400 714 420
rect 714 380 798 400
rect 714 400 798 420
rect 798 380 882 400
rect 798 400 882 420
rect 882 380 966 400
rect 882 400 966 420
rect 966 380 1050 400
rect 966 400 1050 420
rect 1050 380 1134 400
rect 1050 400 1134 420
rect 1134 380 1218 400
rect 1134 400 1218 420
rect 1218 380 1302 400
rect 1218 400 1302 420
rect 1302 380 1386 400
rect 1302 400 1386 420
rect 1386 380 1470 400
rect 1386 400 1470 420
rect 1470 380 1554 400
rect 1470 400 1554 420
rect 1554 380 1596 400
rect 1554 400 1596 420
rect 588 700 630 720
rect 588 720 630 740
rect 630 700 714 720
rect 630 720 714 740
rect 714 700 798 720
rect 714 720 798 740
rect 798 700 882 720
rect 798 720 882 740
rect 882 700 966 720
rect 882 720 966 740
rect 966 700 1050 720
rect 966 720 1050 740
rect 1050 700 1134 720
rect 1050 720 1134 740
rect 1134 700 1218 720
rect 1134 720 1218 740
rect 1218 700 1302 720
rect 1218 720 1302 740
rect 1302 700 1386 720
rect 1302 720 1386 740
rect 1386 700 1470 720
rect 1386 720 1470 740
rect 1470 700 1554 720
rect 1470 720 1554 740
rect 1554 700 1596 720
rect 1554 720 1596 740
<< via1 >>
rect 420 48 462 56
rect 420 56 462 64
rect 420 64 462 72
rect 420 72 462 80
rect 420 80 462 88
rect 420 88 462 96
rect 420 96 462 104
rect 420 104 462 112
rect 462 48 546 56
rect 462 56 546 64
rect 462 64 546 72
rect 462 72 546 80
rect 462 80 546 88
rect 462 88 546 96
rect 462 96 546 104
rect 462 104 546 112
rect 546 48 588 56
rect 546 56 588 64
rect 546 64 588 72
rect 546 72 588 80
rect 546 80 588 88
rect 546 88 588 96
rect 546 96 588 104
rect 546 104 588 112
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1596 368 1638 376
rect 1596 376 1638 384
rect 1596 384 1638 392
rect 1596 392 1638 400
rect 1596 400 1638 408
rect 1596 408 1638 416
rect 1596 416 1638 424
rect 1596 424 1638 432
rect 1638 368 1722 376
rect 1638 376 1722 384
rect 1638 384 1722 392
rect 1638 392 1722 400
rect 1638 400 1722 408
rect 1638 408 1722 416
rect 1638 416 1722 424
rect 1638 424 1722 432
rect 1722 368 1764 376
rect 1722 376 1764 384
rect 1722 384 1764 392
rect 1722 392 1764 400
rect 1722 400 1764 408
rect 1722 408 1764 416
rect 1722 416 1764 424
rect 1722 424 1764 432
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 420 688 462 696
rect 420 696 462 704
rect 420 704 462 712
rect 420 712 462 720
rect 420 720 462 728
rect 420 728 462 736
rect 420 736 462 744
rect 420 744 462 752
rect 462 688 546 696
rect 462 696 546 704
rect 462 704 546 712
rect 462 712 546 720
rect 462 720 546 728
rect 462 728 546 736
rect 462 736 546 744
rect 462 744 546 752
rect 546 688 588 696
rect 546 696 588 704
rect 546 704 588 712
rect 546 712 588 720
rect 546 720 588 728
rect 546 728 588 736
rect 546 736 588 744
rect 546 744 588 752
<< pwell >>
rect -126 -40 2310 840
<< labels >>
flabel metal2 s 210 360 294 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel metal2 s 378 600 630 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel metal1 s -126 360 126 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel metal2 s 1554 40 1806 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2184 800
<< end >>
