magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 1512 480
<< ntap >>
rect -126 120 1638 200
rect -126 200 1638 280
rect -126 280 1638 360
rect -126 360 126 440
rect 1386 360 1638 440
rect -126 440 126 520
rect 1386 440 1638 520
<< metal1 >>
rect -126 120 1638 200
rect -126 200 1638 280
rect -126 280 1638 360
rect -126 360 126 440
rect 1386 360 1638 440
rect -126 440 126 520
rect 1386 440 1638 520
<< ntapc >>
rect 210 200 1218 280
<< nwell >>
rect -210 -124 1722 604
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 1512 480
<< end >>
