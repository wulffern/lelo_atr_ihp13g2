magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 1512 800
<< pdiff >>
rect 546 200 966 280
rect 546 280 966 360
rect 546 360 966 440
rect 546 440 966 520
rect 546 520 966 600
<< ntap >>
rect -126 -40 126 40
rect 1386 -40 1638 40
rect -126 40 126 120
rect 1386 40 1638 120
rect -126 120 126 200
rect 1386 120 1638 200
rect -126 200 126 280
rect 1386 200 1638 280
rect -126 280 126 360
rect 1386 280 1638 360
rect -126 360 126 440
rect 1386 360 1638 440
rect -126 440 126 520
rect 1386 440 1638 520
rect -126 520 126 600
rect 1386 520 1638 600
rect -126 600 126 680
rect 1386 600 1638 680
rect -126 680 126 760
rect 1386 680 1638 760
rect -126 760 126 840
rect 1386 760 1638 840
<< poly >>
rect 210 -14 1302 14
rect 210 146 1302 174
rect 210 306 1302 334
rect 210 466 1302 494
rect 210 626 1302 654
rect 210 786 1302 814
rect 210 280 294 360
rect 1218 280 1302 360
rect 210 360 294 440
rect 1218 360 1302 440
rect 210 440 294 520
rect 1218 440 1302 520
<< metal2 >>
rect 210 360 294 440
rect 378 600 630 680
rect 882 40 1134 120
rect 210 40 294 120
rect 378 40 630 120
rect 882 40 1134 120
rect 210 120 294 200
rect 378 120 630 200
rect 882 120 1134 200
rect 210 200 294 280
rect 378 200 630 280
rect 882 200 1134 280
rect 210 280 294 360
rect 378 280 630 360
rect 882 280 1134 360
rect 210 360 294 440
rect 378 360 630 440
rect 882 360 1134 440
rect 210 440 294 520
rect 378 440 630 520
rect 882 440 1134 520
rect 210 520 294 600
rect 378 520 630 600
rect 882 520 1134 600
rect 210 600 294 680
rect 378 600 630 680
rect 882 600 1134 680
rect 210 680 294 760
rect 378 680 630 760
rect 882 680 1134 760
<< pc >>
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 1232 300 1288 320
rect 1232 320 1288 340
rect 1232 340 1288 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1232 360 1288 380
rect 1232 380 1288 400
rect 1232 400 1288 420
rect 1232 420 1288 440
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 1232 440 1288 460
rect 1232 460 1288 480
rect 1232 480 1288 500
<< metal1 >>
rect -126 -40 126 40
rect 1386 -40 1638 40
rect -126 40 126 120
rect 1386 40 1638 120
rect -126 120 126 200
rect 1386 120 1638 200
rect -126 200 126 280
rect 378 200 966 280
rect 1386 200 1638 280
rect -126 280 126 360
rect 210 280 294 360
rect 1218 280 1302 360
rect 1386 280 1638 360
rect -126 360 126 440
rect -126 360 126 440
rect 210 360 294 440
rect 546 360 1134 440
rect 1218 360 1302 440
rect 1386 360 1638 440
rect -126 440 126 520
rect 210 440 294 520
rect 1218 440 1302 520
rect 1386 440 1638 520
rect -126 520 126 600
rect 378 520 966 600
rect 1386 520 1638 600
rect -126 600 126 680
rect 1386 600 1638 680
rect -126 680 126 760
rect 1386 680 1638 760
rect -126 760 126 840
rect 1386 760 1638 840
<< ntapc >>
rect -42 200 42 280
rect 1470 200 1554 280
rect -42 280 42 360
rect 1470 280 1554 360
rect -42 360 42 440
rect 1470 360 1554 440
rect -42 440 42 520
rect 1470 440 1554 520
rect -42 520 42 600
rect 1470 520 1554 600
<< pdcontact >>
rect 588 220 630 240
rect 588 240 630 260
rect 630 220 714 240
rect 630 240 714 260
rect 714 220 798 240
rect 714 240 798 260
rect 798 220 882 240
rect 798 240 882 260
rect 882 220 924 240
rect 882 240 924 260
rect 588 380 630 400
rect 588 400 630 420
rect 630 380 714 400
rect 630 400 714 420
rect 714 380 798 400
rect 714 400 798 420
rect 798 380 882 400
rect 798 400 882 420
rect 882 380 924 400
rect 882 400 924 420
rect 588 540 630 560
rect 588 560 630 580
rect 630 540 714 560
rect 630 560 714 580
rect 714 540 798 560
rect 714 560 798 580
rect 798 540 882 560
rect 798 560 882 580
rect 882 540 924 560
rect 882 560 924 580
<< via1 >>
rect 420 208 462 216
rect 420 216 462 224
rect 420 224 462 232
rect 420 232 462 240
rect 420 240 462 248
rect 420 248 462 256
rect 420 256 462 264
rect 420 264 462 272
rect 462 208 546 216
rect 462 216 546 224
rect 462 224 546 232
rect 462 232 546 240
rect 462 240 546 248
rect 462 248 546 256
rect 462 256 546 264
rect 462 264 546 272
rect 546 208 588 216
rect 546 216 588 224
rect 546 224 588 232
rect 546 232 588 240
rect 546 240 588 248
rect 546 248 588 256
rect 546 256 588 264
rect 546 264 588 272
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 924 368 966 376
rect 924 376 966 384
rect 924 384 966 392
rect 924 392 966 400
rect 924 400 966 408
rect 924 408 966 416
rect 924 416 966 424
rect 924 424 966 432
rect 966 368 1050 376
rect 966 376 1050 384
rect 966 384 1050 392
rect 966 392 1050 400
rect 966 400 1050 408
rect 966 408 1050 416
rect 966 416 1050 424
rect 966 424 1050 432
rect 1050 368 1092 376
rect 1050 376 1092 384
rect 1050 384 1092 392
rect 1050 392 1092 400
rect 1050 400 1092 408
rect 1050 408 1092 416
rect 1050 416 1092 424
rect 1050 424 1092 432
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 420 528 462 536
rect 420 536 462 544
rect 420 544 462 552
rect 420 552 462 560
rect 420 560 462 568
rect 420 568 462 576
rect 420 576 462 584
rect 420 584 462 592
rect 462 528 546 536
rect 462 536 546 544
rect 462 544 546 552
rect 462 552 546 560
rect 462 560 546 568
rect 462 568 546 576
rect 462 576 546 584
rect 462 584 546 592
rect 546 528 588 536
rect 546 536 588 544
rect 546 544 588 552
rect 546 552 588 560
rect 546 560 588 568
rect 546 568 588 576
rect 546 576 588 584
rect 546 584 588 592
<< nwell >>
rect -210 -124 1722 924
<< labels >>
flabel metal2 s 210 360 294 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel metal2 s 378 600 630 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel metal1 s -126 360 126 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel metal2 s 882 40 1134 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1512 800
<< end >>
