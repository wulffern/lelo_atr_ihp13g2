magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 2688 2560
use LELOATR_PCH_2CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 1344 480
use LELOATR_PCH_2C1F2 xa2 
transform 1 0 0 0 1 480
box 0 480 1344 1280
use LELOATR_PCH_2C5F0 xa3 
transform 1 0 0 0 1 1280
box 0 1280 1344 2080
use LELOATR_PCH_2CTAPTOP xa4 
transform 1 0 0 0 1 2080
box 0 2080 1344 2560
use LELOATR_PCH_2CTAPBOT xb1 
transform 1 0 1344 0 1 0
box 1344 0 2688 480
use LELOATR_PCH_2C1F2 xb2 
transform 1 0 1344 0 1 480
box 1344 480 2688 1280
use LELOATR_PCH_2C5F0 xb3 
transform 1 0 1344 0 1 1280
box 1344 1280 2688 2080
use LELOATR_PCH_2CTAPTOP xb4 
transform 1 0 1344 0 1 2080
box 1344 2080 2688 2560
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 2688 2560
<< end >>
