magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 2184 800
<< pdiff >>
rect 546 200 1638 280
rect 546 280 1638 360
rect 546 360 1638 440
rect 546 440 1638 520
rect 546 520 1638 600
<< ntap >>
rect -126 -40 126 40
rect 2058 -40 2310 40
rect -126 40 126 120
rect 2058 40 2310 120
rect -126 120 126 200
rect 2058 120 2310 200
rect -126 200 126 280
rect 2058 200 2310 280
rect -126 280 126 360
rect 2058 280 2310 360
rect -126 360 126 440
rect 2058 360 2310 440
rect -126 440 126 520
rect 2058 440 2310 520
rect -126 520 126 600
rect 2058 520 2310 600
rect -126 600 126 680
rect 2058 600 2310 680
rect -126 680 126 760
rect 2058 680 2310 760
rect -126 760 126 840
rect 2058 760 2310 840
<< poly >>
rect 210 -14 1974 14
rect 210 146 1974 174
rect 210 306 1974 334
rect 210 466 1974 494
rect 210 626 1974 654
rect 210 786 1974 814
rect 210 280 294 360
rect 1890 280 1974 360
rect 210 360 294 440
rect 1890 360 1974 440
rect 210 440 294 520
rect 1890 440 1974 520
<< metal2 >>
rect 210 360 294 440
rect 378 600 630 680
rect 1554 40 1806 120
rect 210 40 294 120
rect 378 40 630 120
rect 1554 40 1806 120
rect 210 120 294 200
rect 378 120 630 200
rect 1554 120 1806 200
rect 210 200 294 280
rect 378 200 630 280
rect 1554 200 1806 280
rect 210 280 294 360
rect 378 280 630 360
rect 1554 280 1806 360
rect 210 360 294 440
rect 378 360 630 440
rect 1554 360 1806 440
rect 210 440 294 520
rect 378 440 630 520
rect 1554 440 1806 520
rect 210 520 294 600
rect 378 520 630 600
rect 1554 520 1806 600
rect 210 600 294 680
rect 378 600 630 680
rect 1554 600 1806 680
rect 210 680 294 760
rect 378 680 630 760
rect 1554 680 1806 760
<< pc >>
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 1904 300 1960 320
rect 1904 320 1960 340
rect 1904 340 1960 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1904 360 1960 380
rect 1904 380 1960 400
rect 1904 400 1960 420
rect 1904 420 1960 440
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 1904 440 1960 460
rect 1904 460 1960 480
rect 1904 480 1960 500
<< metal1 >>
rect -126 -40 126 40
rect 2058 -40 2310 40
rect -126 40 126 120
rect 2058 40 2310 120
rect -126 120 126 200
rect 2058 120 2310 200
rect -126 200 126 280
rect 378 200 1638 280
rect 2058 200 2310 280
rect -126 280 126 360
rect 210 280 294 360
rect 1890 280 1974 360
rect 2058 280 2310 360
rect -126 360 126 440
rect -126 360 126 440
rect 210 360 294 440
rect 546 360 1806 440
rect 1890 360 1974 440
rect 2058 360 2310 440
rect -126 440 126 520
rect 210 440 294 520
rect 1890 440 1974 520
rect 2058 440 2310 520
rect -126 520 126 600
rect 378 520 1638 600
rect 2058 520 2310 600
rect -126 600 126 680
rect 2058 600 2310 680
rect -126 680 126 760
rect 2058 680 2310 760
rect -126 760 126 840
rect 2058 760 2310 840
<< ntapc >>
rect -42 200 42 280
rect 2142 200 2226 280
rect -42 280 42 360
rect 2142 280 2226 360
rect -42 360 42 440
rect 2142 360 2226 440
rect -42 440 42 520
rect 2142 440 2226 520
rect -42 520 42 600
rect 2142 520 2226 600
<< pdcontact >>
rect 588 220 630 240
rect 588 240 630 260
rect 630 220 714 240
rect 630 240 714 260
rect 714 220 798 240
rect 714 240 798 260
rect 798 220 882 240
rect 798 240 882 260
rect 882 220 966 240
rect 882 240 966 260
rect 966 220 1050 240
rect 966 240 1050 260
rect 1050 220 1134 240
rect 1050 240 1134 260
rect 1134 220 1218 240
rect 1134 240 1218 260
rect 1218 220 1302 240
rect 1218 240 1302 260
rect 1302 220 1386 240
rect 1302 240 1386 260
rect 1386 220 1470 240
rect 1386 240 1470 260
rect 1470 220 1554 240
rect 1470 240 1554 260
rect 1554 220 1596 240
rect 1554 240 1596 260
rect 588 380 630 400
rect 588 400 630 420
rect 630 380 714 400
rect 630 400 714 420
rect 714 380 798 400
rect 714 400 798 420
rect 798 380 882 400
rect 798 400 882 420
rect 882 380 966 400
rect 882 400 966 420
rect 966 380 1050 400
rect 966 400 1050 420
rect 1050 380 1134 400
rect 1050 400 1134 420
rect 1134 380 1218 400
rect 1134 400 1218 420
rect 1218 380 1302 400
rect 1218 400 1302 420
rect 1302 380 1386 400
rect 1302 400 1386 420
rect 1386 380 1470 400
rect 1386 400 1470 420
rect 1470 380 1554 400
rect 1470 400 1554 420
rect 1554 380 1596 400
rect 1554 400 1596 420
rect 588 540 630 560
rect 588 560 630 580
rect 630 540 714 560
rect 630 560 714 580
rect 714 540 798 560
rect 714 560 798 580
rect 798 540 882 560
rect 798 560 882 580
rect 882 540 966 560
rect 882 560 966 580
rect 966 540 1050 560
rect 966 560 1050 580
rect 1050 540 1134 560
rect 1050 560 1134 580
rect 1134 540 1218 560
rect 1134 560 1218 580
rect 1218 540 1302 560
rect 1218 560 1302 580
rect 1302 540 1386 560
rect 1302 560 1386 580
rect 1386 540 1470 560
rect 1386 560 1470 580
rect 1470 540 1554 560
rect 1470 560 1554 580
rect 1554 540 1596 560
rect 1554 560 1596 580
<< via1 >>
rect 420 208 462 216
rect 420 216 462 224
rect 420 224 462 232
rect 420 232 462 240
rect 420 240 462 248
rect 420 248 462 256
rect 420 256 462 264
rect 420 264 462 272
rect 462 208 546 216
rect 462 216 546 224
rect 462 224 546 232
rect 462 232 546 240
rect 462 240 546 248
rect 462 248 546 256
rect 462 256 546 264
rect 462 264 546 272
rect 546 208 588 216
rect 546 216 588 224
rect 546 224 588 232
rect 546 232 588 240
rect 546 240 588 248
rect 546 248 588 256
rect 546 256 588 264
rect 546 264 588 272
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1596 368 1638 376
rect 1596 376 1638 384
rect 1596 384 1638 392
rect 1596 392 1638 400
rect 1596 400 1638 408
rect 1596 408 1638 416
rect 1596 416 1638 424
rect 1596 424 1638 432
rect 1638 368 1722 376
rect 1638 376 1722 384
rect 1638 384 1722 392
rect 1638 392 1722 400
rect 1638 400 1722 408
rect 1638 408 1722 416
rect 1638 416 1722 424
rect 1638 424 1722 432
rect 1722 368 1764 376
rect 1722 376 1764 384
rect 1722 384 1764 392
rect 1722 392 1764 400
rect 1722 400 1764 408
rect 1722 408 1764 416
rect 1722 416 1764 424
rect 1722 424 1764 432
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 420 528 462 536
rect 420 536 462 544
rect 420 544 462 552
rect 420 552 462 560
rect 420 560 462 568
rect 420 568 462 576
rect 420 576 462 584
rect 420 584 462 592
rect 462 528 546 536
rect 462 536 546 544
rect 462 544 546 552
rect 462 552 546 560
rect 462 560 546 568
rect 462 568 546 576
rect 462 576 546 584
rect 462 584 546 592
rect 546 528 588 536
rect 546 536 588 544
rect 546 544 588 552
rect 546 552 588 560
rect 546 560 588 568
rect 546 568 588 576
rect 546 576 588 584
rect 546 584 588 592
<< nwell >>
rect -210 -124 2394 924
<< labels >>
flabel metal2 s 210 360 294 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel metal2 s 378 600 630 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel metal1 s -126 360 126 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel metal2 s 1554 40 1806 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 2184 800
<< end >>
