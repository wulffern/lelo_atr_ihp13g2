magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 1344 800
<< pdiff >>
rect 546 40 798 120
rect 546 120 798 200
rect 546 200 798 280
rect 546 280 798 360
rect 546 360 798 440
rect 546 440 798 520
rect 546 520 798 600
rect 546 600 798 680
rect 546 680 798 760
<< ptap >>
rect -126 -40 126 40
rect 1218 -40 1470 40
rect -126 40 126 120
rect 1218 40 1470 120
rect -126 120 126 200
rect 1218 120 1470 200
rect -126 200 126 280
rect 1218 200 1470 280
rect -126 280 126 360
rect 1218 280 1470 360
rect -126 360 126 440
rect 1218 360 1470 440
rect -126 440 126 520
rect 1218 440 1470 520
rect -126 520 126 600
rect 1218 520 1470 600
rect -126 600 126 680
rect 1218 600 1470 680
rect -126 680 126 760
rect 1218 680 1470 760
rect -126 760 126 840
rect 1218 760 1470 840
<< poly >>
rect 210 140 1134 340
rect 210 460 1134 660
rect 210 -14 1134 14
rect 210 200 294 280
rect 1050 200 1134 280
rect 210 280 294 360
rect 1050 280 1134 360
rect 210 360 294 440
rect 1050 360 1134 440
rect 210 440 294 520
rect 1050 440 1134 520
rect 210 520 294 600
rect 1050 520 1134 600
rect 210 786 1134 814
<< metal2 >>
rect 210 360 294 440
rect 378 600 630 680
rect 714 40 966 120
rect 210 40 294 120
rect 378 40 630 120
rect 714 40 966 120
rect 210 120 294 200
rect 378 120 630 200
rect 714 120 966 200
rect 210 200 294 280
rect 378 200 630 280
rect 714 200 966 280
rect 210 280 294 360
rect 378 280 630 360
rect 714 280 966 360
rect 210 360 294 440
rect 378 360 630 440
rect 714 360 966 440
rect 210 440 294 520
rect 378 440 630 520
rect 714 440 966 520
rect 210 520 294 600
rect 378 520 630 600
rect 714 520 966 600
rect 210 600 294 680
rect 378 600 630 680
rect 714 600 966 680
rect 210 680 294 760
rect 378 680 630 760
rect 714 680 966 760
<< pc >>
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 1064 300 1120 320
rect 1064 320 1120 340
rect 1064 340 1120 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1064 360 1120 380
rect 1064 380 1120 400
rect 1064 400 1120 420
rect 1064 420 1120 440
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 1064 440 1120 460
rect 1064 460 1120 480
rect 1064 480 1120 500
<< metal1 >>
rect -126 -40 126 40
rect 1218 -40 1470 40
rect -126 40 126 120
rect 378 40 798 120
rect 1218 40 1470 120
rect -126 120 126 200
rect 1218 120 1470 200
rect -126 200 126 280
rect 1218 200 1470 280
rect -126 280 126 360
rect 210 280 294 360
rect 1050 280 1134 360
rect 1218 280 1470 360
rect -126 360 126 440
rect -126 360 126 440
rect 210 360 294 440
rect 546 360 966 440
rect 1050 360 1134 440
rect 1218 360 1470 440
rect -126 440 126 520
rect 210 440 294 520
rect 1050 440 1134 520
rect 1218 440 1470 520
rect -126 520 126 600
rect 1218 520 1470 600
rect -126 600 126 680
rect 1218 600 1470 680
rect -126 680 126 760
rect 378 680 798 760
rect 1218 680 1470 760
rect -126 760 126 840
rect 1218 760 1470 840
<< ptapc >>
rect -42 200 42 280
rect 1302 200 1386 280
rect -42 280 42 360
rect 1302 280 1386 360
rect -42 360 42 440
rect 1302 360 1386 440
rect -42 440 42 520
rect 1302 440 1386 520
rect -42 520 42 600
rect 1302 520 1386 600
<< ndcontact >>
rect 588 60 630 80
rect 588 80 630 100
rect 630 60 714 80
rect 630 80 714 100
rect 714 60 756 80
rect 714 80 756 100
rect 588 380 630 400
rect 588 400 630 420
rect 630 380 714 400
rect 630 400 714 420
rect 714 380 756 400
rect 714 400 756 420
rect 588 700 630 720
rect 588 720 630 740
rect 630 700 714 720
rect 630 720 714 740
rect 714 700 756 720
rect 714 720 756 740
<< via1 >>
rect 420 48 462 56
rect 420 56 462 64
rect 420 64 462 72
rect 420 72 462 80
rect 420 80 462 88
rect 420 88 462 96
rect 420 96 462 104
rect 420 104 462 112
rect 462 48 546 56
rect 462 56 546 64
rect 462 64 546 72
rect 462 72 546 80
rect 462 80 546 88
rect 462 88 546 96
rect 462 96 546 104
rect 462 104 546 112
rect 546 48 588 56
rect 546 56 588 64
rect 546 64 588 72
rect 546 72 588 80
rect 546 80 588 88
rect 546 88 588 96
rect 546 96 588 104
rect 546 104 588 112
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 756 368 798 376
rect 756 376 798 384
rect 756 384 798 392
rect 756 392 798 400
rect 756 400 798 408
rect 756 408 798 416
rect 756 416 798 424
rect 756 424 798 432
rect 798 368 882 376
rect 798 376 882 384
rect 798 384 882 392
rect 798 392 882 400
rect 798 400 882 408
rect 798 408 882 416
rect 798 416 882 424
rect 798 424 882 432
rect 882 368 924 376
rect 882 376 924 384
rect 882 384 924 392
rect 882 392 924 400
rect 882 400 924 408
rect 882 408 924 416
rect 882 416 924 424
rect 882 424 924 432
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 420 688 462 696
rect 420 696 462 704
rect 420 704 462 712
rect 420 712 462 720
rect 420 720 462 728
rect 420 728 462 736
rect 420 736 462 744
rect 420 744 462 752
rect 462 688 546 696
rect 462 696 546 704
rect 462 704 546 712
rect 462 712 546 720
rect 462 720 546 728
rect 462 728 546 736
rect 462 736 546 744
rect 462 744 546 752
rect 546 688 588 696
rect 546 696 588 704
rect 546 704 588 712
rect 546 712 588 720
rect 546 720 588 728
rect 546 728 588 736
rect 546 736 588 744
rect 546 744 588 752
<< pwell >>
rect -126 -40 1470 840
<< labels >>
flabel metal2 s 210 360 294 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel metal2 s 378 600 630 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel metal1 s -126 360 126 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel metal2 s 714 40 966 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1344 800
<< end >>
