magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 1512 480
<< ptap >>
rect -126 -40 126 40
rect 1386 -40 1638 40
rect -126 40 126 120
rect 1386 40 1638 120
rect -126 120 1638 200
rect -126 200 1638 280
rect -126 280 1638 360
<< metal1 >>
rect -126 -40 126 40
rect 1386 -40 1638 40
rect -126 40 126 120
rect 1386 40 1638 120
rect -126 120 1638 200
rect -126 200 1638 280
rect -126 280 1638 360
<< ptapc >>
rect 210 200 1302 280
<< pwell >>
rect -126 -40 1638 520
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 1512 480
<< end >>
