magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 1848 800
<< pdiff >>
rect 546 40 1302 120
rect 546 120 1302 200
rect 546 200 1302 280
rect 546 280 1302 360
rect 546 360 1302 440
rect 546 440 1302 520
rect 546 520 1302 600
rect 546 600 1302 680
rect 546 680 1302 760
<< ptap >>
rect -126 -40 126 40
rect 1722 -40 1974 40
rect -126 40 126 120
rect 1722 40 1974 120
rect -126 120 126 200
rect 1722 120 1974 200
rect -126 200 126 280
rect 1722 200 1974 280
rect -126 280 126 360
rect 1722 280 1974 360
rect -126 360 126 440
rect 1722 360 1974 440
rect -126 440 126 520
rect 1722 440 1974 520
rect -126 520 126 600
rect 1722 520 1974 600
rect -126 600 126 680
rect 1722 600 1974 680
rect -126 680 126 760
rect 1722 680 1974 760
rect -126 760 126 840
rect 1722 760 1974 840
<< poly >>
rect 210 140 1638 340
rect 210 460 1638 660
rect 210 -14 1638 14
rect 210 200 294 280
rect 1554 200 1638 280
rect 210 280 294 360
rect 1554 280 1638 360
rect 210 360 294 440
rect 1554 360 1638 440
rect 210 440 294 520
rect 1554 440 1638 520
rect 210 520 294 600
rect 1554 520 1638 600
rect 210 786 1638 814
<< metal2 >>
rect 210 360 294 440
rect 378 600 630 680
rect 1218 40 1470 120
rect 210 40 294 120
rect 378 40 630 120
rect 1218 40 1470 120
rect 210 120 294 200
rect 378 120 630 200
rect 1218 120 1470 200
rect 210 200 294 280
rect 378 200 630 280
rect 1218 200 1470 280
rect 210 280 294 360
rect 378 280 630 360
rect 1218 280 1470 360
rect 210 360 294 440
rect 378 360 630 440
rect 1218 360 1470 440
rect 210 440 294 520
rect 378 440 630 520
rect 1218 440 1470 520
rect 210 520 294 600
rect 378 520 630 600
rect 1218 520 1470 600
rect 210 600 294 680
rect 378 600 630 680
rect 1218 600 1470 680
rect 210 680 294 760
rect 378 680 630 760
rect 1218 680 1470 760
<< pc >>
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 1568 300 1624 320
rect 1568 320 1624 340
rect 1568 340 1624 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1568 360 1624 380
rect 1568 380 1624 400
rect 1568 400 1624 420
rect 1568 420 1624 440
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 1568 440 1624 460
rect 1568 460 1624 480
rect 1568 480 1624 500
<< metal1 >>
rect -126 -40 126 40
rect 1722 -40 1974 40
rect -126 40 126 120
rect 378 40 1302 120
rect 1722 40 1974 120
rect -126 120 126 200
rect 1722 120 1974 200
rect -126 200 126 280
rect 1722 200 1974 280
rect -126 280 126 360
rect 210 280 294 360
rect 1554 280 1638 360
rect 1722 280 1974 360
rect -126 360 126 440
rect -126 360 126 440
rect 210 360 294 440
rect 546 360 1470 440
rect 1554 360 1638 440
rect 1722 360 1974 440
rect -126 440 126 520
rect 210 440 294 520
rect 1554 440 1638 520
rect 1722 440 1974 520
rect -126 520 126 600
rect 1722 520 1974 600
rect -126 600 126 680
rect 1722 600 1974 680
rect -126 680 126 760
rect 378 680 1302 760
rect 1722 680 1974 760
rect -126 760 126 840
rect 1722 760 1974 840
<< ptapc >>
rect -42 200 42 280
rect 1806 200 1890 280
rect -42 280 42 360
rect 1806 280 1890 360
rect -42 360 42 440
rect 1806 360 1890 440
rect -42 440 42 520
rect 1806 440 1890 520
rect -42 520 42 600
rect 1806 520 1890 600
<< ndcontact >>
rect 588 60 630 80
rect 588 80 630 100
rect 630 60 714 80
rect 630 80 714 100
rect 714 60 798 80
rect 714 80 798 100
rect 798 60 882 80
rect 798 80 882 100
rect 882 60 966 80
rect 882 80 966 100
rect 966 60 1050 80
rect 966 80 1050 100
rect 1050 60 1134 80
rect 1050 80 1134 100
rect 1134 60 1218 80
rect 1134 80 1218 100
rect 1218 60 1260 80
rect 1218 80 1260 100
rect 588 380 630 400
rect 588 400 630 420
rect 630 380 714 400
rect 630 400 714 420
rect 714 380 798 400
rect 714 400 798 420
rect 798 380 882 400
rect 798 400 882 420
rect 882 380 966 400
rect 882 400 966 420
rect 966 380 1050 400
rect 966 400 1050 420
rect 1050 380 1134 400
rect 1050 400 1134 420
rect 1134 380 1218 400
rect 1134 400 1218 420
rect 1218 380 1260 400
rect 1218 400 1260 420
rect 588 700 630 720
rect 588 720 630 740
rect 630 700 714 720
rect 630 720 714 740
rect 714 700 798 720
rect 714 720 798 740
rect 798 700 882 720
rect 798 720 882 740
rect 882 700 966 720
rect 882 720 966 740
rect 966 700 1050 720
rect 966 720 1050 740
rect 1050 700 1134 720
rect 1050 720 1134 740
rect 1134 700 1218 720
rect 1134 720 1218 740
rect 1218 700 1260 720
rect 1218 720 1260 740
<< via1 >>
rect 420 48 462 56
rect 420 56 462 64
rect 420 64 462 72
rect 420 72 462 80
rect 420 80 462 88
rect 420 88 462 96
rect 420 96 462 104
rect 420 104 462 112
rect 462 48 546 56
rect 462 56 546 64
rect 462 64 546 72
rect 462 72 546 80
rect 462 80 546 88
rect 462 88 546 96
rect 462 96 546 104
rect 462 104 546 112
rect 546 48 588 56
rect 546 56 588 64
rect 546 64 588 72
rect 546 72 588 80
rect 546 80 588 88
rect 546 88 588 96
rect 546 96 588 104
rect 546 104 588 112
rect 224 300 280 320
rect 224 320 280 340
rect 224 340 280 360
rect 224 360 280 380
rect 224 380 280 400
rect 224 400 280 420
rect 224 420 280 440
rect 1260 368 1302 376
rect 1260 376 1302 384
rect 1260 384 1302 392
rect 1260 392 1302 400
rect 1260 400 1302 408
rect 1260 408 1302 416
rect 1260 416 1302 424
rect 1260 424 1302 432
rect 1302 368 1386 376
rect 1302 376 1386 384
rect 1302 384 1386 392
rect 1302 392 1386 400
rect 1302 400 1386 408
rect 1302 408 1386 416
rect 1302 416 1386 424
rect 1302 424 1386 432
rect 1386 368 1428 376
rect 1386 376 1428 384
rect 1386 384 1428 392
rect 1386 392 1428 400
rect 1386 400 1428 408
rect 1386 408 1428 416
rect 1386 416 1428 424
rect 1386 424 1428 432
rect 224 440 280 460
rect 224 460 280 480
rect 224 480 280 500
rect 420 688 462 696
rect 420 696 462 704
rect 420 704 462 712
rect 420 712 462 720
rect 420 720 462 728
rect 420 728 462 736
rect 420 736 462 744
rect 420 744 462 752
rect 462 688 546 696
rect 462 696 546 704
rect 462 704 546 712
rect 462 712 546 720
rect 462 720 546 728
rect 462 728 546 736
rect 462 736 546 744
rect 462 744 546 752
rect 546 688 588 696
rect 546 696 588 704
rect 546 704 588 712
rect 546 712 588 720
rect 546 720 588 728
rect 546 728 588 736
rect 546 736 588 744
rect 546 744 588 752
<< pwell >>
rect -126 -40 1974 840
<< labels >>
flabel metal2 s 210 360 294 440 0 FreeSans 400 0 0 0 G
port 2 nsew signal bidirectional
flabel metal2 s 378 600 630 680 0 FreeSans 400 0 0 0 S
port 3 nsew signal bidirectional
flabel metal1 s -126 360 126 440 0 FreeSans 400 0 0 0 B
port 4 nsew signal bidirectional
flabel metal2 s 1218 40 1470 120 0 FreeSans 400 0 0 0 D
port 1 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 1848 800
<< end >>
