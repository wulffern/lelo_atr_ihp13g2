magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741993200
<< checkpaint >>
rect 0 0 4368 2560
use LELOATR_NCH_12CTAPBOT xa1 
transform 1 0 0 0 1 0
box 0 0 2184 480
use LELOATR_NCH_12C1F2 xa2 
transform 1 0 0 0 1 480
box 0 480 2184 1280
use LELOATR_NCH_12C5F0 xa3 
transform 1 0 0 0 1 1280
box 0 1280 2184 2080
use LELOATR_NCH_12CTAPTOP xa4 
transform 1 0 0 0 1 2080
box 0 2080 2184 2560
use LELOATR_NCH_12CTAPBOT xb1 
transform 1 0 2184 0 1 0
box 2184 0 4368 480
use LELOATR_NCH_12C1F2 xb2 
transform 1 0 2184 0 1 480
box 2184 480 4368 1280
use LELOATR_NCH_12C5F0 xb3 
transform 1 0 2184 0 1 1280
box 2184 1280 4368 2080
use LELOATR_NCH_12CTAPTOP xb4 
transform 1 0 2184 0 1 2080
box 2184 2080 4368 2560
<< labels >>
<< properties >>
string FIXED_BBOX 0 0 4368 2560
<< end >>
